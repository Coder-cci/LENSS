Begin3
Language:    SV, 850, Swedish
Title:       shext
Description: Share Extender
Keywords:    delning ut�kning
End
