Begin3
Language:    SV, 850, Swedish
Title:       SHSUFDRV
Description: SHSUFDRV �r en drivrutin f�r diskett- och h�rddiskavbildningar. SHSURDRV kopierar avbildningen till RAM och/eller skapar RAM-enheter.
Keywords:    drivrutin, diskett, avbildningar, h�rddisk, ramdisk
End
