Begin3
Language:    SV, 850, Swedish
Title:       Crynwr
Description: En samling av fria paketdrivrutiner fr�n f�retaget Crynwr
Keywords:    paket
End
