Begin3
Language:    SV, 850, Swedish
Description: Flyttar filer h�rifr�n till dit
Keywords:    freedos, move, flytta
End
