Begin3
Language:    SV, 850, Swedish
Title:       lzop
Description: En komprimerare i stil med gzip, som v�rdes�tter hastighet �ver kompressionsgrad
Keywords:    lzop, kompression
End
