Begin3
Language:    SV, 850, Swedish
Title:       NewSNUZ
Description: Usenet-l�sare (NNTP) baserad p� WatTCP
Keywords:    nntp,usenet
End
