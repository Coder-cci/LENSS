Begin3
Language:    SV, 850, Swedish
Title:       choice
Description: Presentera ett alternativ f�r anv�ndaren och v�nta p� en tangent (anv�nder kitte ist�llet f�r cats)
Keywords:    freedos
End
