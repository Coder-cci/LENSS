Begin3
Language:    SV, 850, Swedish
Title:       KRaptor
Description: Kraptor �r ett Raptor-liknande spel med �ppen k�llkod, komplett med flera banor.
Keywords:    raptor, spel, skjutspel
End
