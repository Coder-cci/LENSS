Begin3
Language:    SV, 850, Swedish
Title:       Mirror
Description: Spelar in information om disken f�r eventuellt data�terst�llning.
Keywords:    freedos
End
