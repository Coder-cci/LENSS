Begin3
Language:    SV, 850, Swedish
Description: FreeDOS installationsprogram - min programvara f�r paketlistredigering
Summary:     FDIMPLES �r paketlistredigeraren f�r det avancerade l�get i FreeDOS installationsprogrammet (FDI). Den kan k�ra som ett separat program som ett mer anv�ndarv�nligt gr�nssnitt till pakethanterarverktyget FDINST som k�r p� kommandoraden.
Keywords:    dos 16-bitars, asm, pascal
End
