Begin3
Language:    SV, 850, Swedish
Title:       which
Description: which �r ett verktyg fr�n UNIX-v�rlden som l�ter anv�ndare hitta k�rbara filer i katalogerna listade i milj�variabeln PATH. Fullt st�d f�r jokertecken, relativa s�kv�gare, valfria fildetaljer (storlek, datum). Anv�ndardefinierbara program�ndelser, kodsides-korreka tids-/datumformatering. Nytt DOS sitchar-st�d.
Keywords:    DOS, ut�kning, fil, verktyg, hitta, PATH
End
