Begin3
Language:    SV, 850, Swedish
Title:       hangman
Description: Flerspr�kig h�nga gubben
Keywords:    h�nga gubbe
End
