Begin3
Language:    SV, 850, Swedish
Title:       XCopy
Description: Kopierar filer och katalogstr�d.
Keywords:    freedos, kopiera, xcopy, kitten
End
