Begin3
Language:    SV, 850, Swedish
Description: Allm�nna underh�llsverktyg f�r FreeDOS-paket
Summary:     Verktyg f�r att skapa och visa information om installerade paket f�r FreeDOS. S� sm�ningom kan verktyg f�r att omplacera, ta bort och utf�ra annat allm�nt paketunderh�ll komma att l�ggas till.
Keywords:    dos 16-bitars, asm, pascal
End
