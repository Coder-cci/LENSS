Begin3
Language:    SV, 850, Swedish
Title:       UHDD
Description: UHDD �r en cachande drivrutin f�r upp till 10 BIOS h�rddiskar/SSD p� upp till 4 UltraDMA-styrkort. Det kommer ocks� att tillhandah�lla cachning f�r diskar som hanteras av UDVD2 om det l�ses in efter UHDD.
Keywords:    cache, disk, dma, drivrutin, ide, sata, ultradma
End
