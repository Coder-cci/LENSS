Begin3
Language:    SV, 850, Swedish
Title:       REPLACE
Description: Ers�tter filer i destinationskatalogen med filer fr�n k�llkatalogen som har samma namn.
Keywords:    kopiera, ers�tt
End
