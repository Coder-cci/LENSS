Begin3
Language:    SV, 850, Swedish
Title:       Eliza
Description: En av de tidigaste datorbaserade AI-tjattrobotarna
End
