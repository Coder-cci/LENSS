Begin3
Language:    SV, 850, Swedish
Title:       Spool
Description: Spolar filutskrifter i bakgrunden. Detta kr�ver inte anv�ndning av PRINT-kommandot.
Keywords:    skriv ut, spooler
End
