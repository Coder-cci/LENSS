Begin3
Language:    SV, 850, Swedish
Title:       Wing
Description: Ett galaga-liknanan rymdskjutspel.
Keywords:    galaga
End
