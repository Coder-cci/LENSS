Begin3
Language:    SV, 850, Swedish
Title:       TOUCH
Description: S�tter datum- och tidst�mplar p� filer likt touch i *nix
Keywords:    touch, tidsst�mpel, unix
End
