Begin3
Language:    SV, 850, Swedish
Title:       GNU sed
Description: GNU sed �r en GNU-implementation av POSIX str�mredigerarer `sed'.
Keywords:    sed
End
