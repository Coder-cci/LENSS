Begin3
Language:    SV, 850, Swedish
Title:       File Slicer
Description: Ett enkelt DOS-arkivverktyg som ocks� kan dela och �terkombinera filer. (UPX-komprimerat)
Summary:     Ett enkelt arkivverktyg (inte ett filkompressionsprogram) f�r att kategoriser och dela stora filer och kataloger �ver mindre media. Det kr�ver en 8086 med EGA-grafik eller b�ttr. (UPX-komprimerat)
Keywords:    dos 16-bitars filarkiv dela upp dela
End
