Begin3
Language:    SV, 850, Swedish
Description: 32-bitars DPI DOS extender designad f�r DJGPP.
End
