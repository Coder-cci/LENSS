# Translation by Martin Str�mberg <ams@ludd.luth.se>.
0.0:Visar alla rader i en fil som inneh�ller en viss str�ng
0.1:R�kna antalet g�nger str�ngen f�rekommer
0.2:Hantera versaler och gemener som lika
0.3:Numrera de visade raderna med start fr�n 1
0.4:Visa raderna som inte inneh�ller str�ngen
1.0:fil
1.1:str�ng
2.0:Kan inte �ppna filen
2.1:Ingen s�dan fil
2.2:Kan inte byta till katalog
