Begin3
Language:    SV, 850, Swedish
Title:       GCDROM
Description: SATA inbyggd IDE CD/DVD-ROM-drivrutin f�r DOS (ocks� k�nd som 'ODD DOS-drivrutin') med st�d f�r alla SATA inbyggda IDE-styrkort s� som Intel ICH6/ICH7/ICH8, Jmicron 363/368, Nvidia CK804 MCP55/MCP51 etc. (byggt fr�n XCDROM med �ndrat namn)
Keywords:    CD-ROM drivrutin, SATA, drivrutin
End
