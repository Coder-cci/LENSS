Begin3
Language:    SV, 850, Swedish
Title:       BladeEnc
Description: Blade's MP3 Encoder genererar MP3-filer fr�n WAV/AIFF/RAW-data
Keywords:    mp3, kodare
End
