Begin3
Language:    SV, 850, Swedish
Title:       OpenCubic Player
Description: OpenCubic Player �r en musikspelare f�r m�nga format (mp3,wav,mid...)
Keywords:    spelare
End
