# Hj�lpmeddelande

0.0:Anv�ndning: MD5SUM [/TBV] [/C [fil]] | [fil...]
0.1:Genererar eller kontrollerar MD5 kontrollsummor
0.2:    /C           kontrollera kontrollsumma (standard �r generera)
0.3:    /[-]V        (in-)aktivera utf�rligt l�ge (standard �r av)
0.4:    /[-]L        (in-)aktivera LFN-anv�ndning (standard �r aktivt)
0.5:    /[-]R[num]   (in-)aktivera rekursion (standard �r av), num �r
0.6:                 ett tal mellan 1-9 som begr�nsar rekursionen (standard=4)
0.7:    /[-]S        samma som /[-]R=]
0.8:    /T           l�ser filer i textl�ge
0.9:    /B           l�ser filer i bin�rt l�ge (standard; �sidos�tts av /T)
0.10:    /M[:|=]l�ge  v�ljer l�ge f�r kontrollsumma (SHA eller MD5)
0.11:Indatan till /C ska vara en lista av kontrollsummor och filnamn som skrivits
0.12:ut p� standard ut av detta program n�r det genererat kontrollsummor.
0.13:Argumentet till /M ska vara ett l�ge, vilket kan vara SHA, CRC32
0.14:SHA256 eller MD5, beroende p� hur MD5SUM kompilerats.

# Diverse andra meddelanden

1.0:Ogiltig flagga in
1.1:File existerar inte
1.2:l�sfel p� standard in
1.3:fel vid l�sning
1.4:ok�nd rad
1.5:kan inte �ppna
1.6:MISSLYCKADES
1.7:kontroll misslyckades f�r
1.8:av
1.9:fil(er) misslyckades i kontroll
1.10:inga filer kontrollerade
1.11:Filen �r en underkatalog
1.12:Varning: LFN st�ds ej
1.13:Flagga saknar argument
1.14:Ogiltigt l�ge f�r kontrollsumma
1.15:Katalog existerar ej
1.16:Kunde inte h�mta den aktuella katalogen
