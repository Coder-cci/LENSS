Begin3
Language:    SV, 850, Swedish
Title:       rsync
Description: rsync �r en verktygsprogramvara som synkroniserar filer och kataloger fr�n en plats til en annan medan det minimerar data�verf�ring genom deltakodning n�r s� �r l�mpligt. Denna rsync-portering �r n�dv�ndigtvis en delm�ngd av den fulla rsync, delvis p� grund av minnebegr�nsningar och delvis p� grund av egenheter hos DOS. Huvudskillnaderna �r: Endast f�r klient; inget st�d f�r rsh eller ssh; filnamn p� servern m�ste vara i DOS-format; fildata komprimeras inte.
Keywords:    rsync
End
