Begin3
Language:    SV, 850, Swedish
Title:       picoTCP
Description: picoTCP-n�tverksstack (bibliotek och konfigurationsverktyg)
End
