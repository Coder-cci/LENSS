Begin3
Language:    SV, 850, Swedish
Title:       FDNPKG
Description: N�tverksbaserad pakethanterare
Keywords:    fdnpkg,uppdatering,paket
End
