Begin3
Language:    SV, 850, Swedish
Title:       Vitetris
Description: En terminal-baserad Tetris-klon.
End
