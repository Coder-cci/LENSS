Begin3
Language:    SV, 850, Swedish
Title:       HEAD
Description: Visar en del av en fil
Keywords:    head
End
