Begin3
Language:    SV, 850, Swedish
Title:       COMP
Description: J�mf�r filer och visa deras skillnader
Keywords:    j�mf�r, comp, filj�mf�relse
End
