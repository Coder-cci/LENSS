Begin3
Language:    SV, 850, Swedish
Title:       sudoku86
Description: Ett 16-bitars Sudoku-spel f�r DOS och 8086/8088 CPU:er
Keywords:    sudoku,spel
End
