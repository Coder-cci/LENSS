Begin3
Language:    SV, 850, Swedish
Title:       CHKDSK
Description: Kontrollera disken efter fel.
Keywords:    kontrollera diskfel
End
