Begin3
Language:    SV, 850, Swedish
Title:       NTFS
Description: M�jligg�r �tkomst av NTFS-partitioner
Keywords:    ntfs, partition, fil, �tkomst
End
