Begin3
Language:    SV, 850, Swedish
Description: DOSSHELL grafiskt anv�ndargr�nssnit implementerat f�r FreeDOS
End
