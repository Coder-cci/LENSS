Begin3
Language:    SV, 850, Swedish
Title:       NetHack
Description: Ett spel f�r en spelare som utforskar en grotta.
End
