Begin3
Language:    SV, 850, Swedish
Title:       NLSFunc
Description: NLSFUNC l�gger till NLS-funktionalitet (Nationellt spr�kst�d)
Keywords:    freedos, nls, country, visa, l�ge
End
