Begin3
Language:    SV, 850, Swedish
Title:       fdxms
Description: Ers�ttnings-drivrutin f�r XMS f�r '386-system eller b�ttre
Keywords:    freedos, xms, himem
End
