Begin3
Language:    SV, 850, Swedish
Title:       M2WAT
Description: Verktyg f�r att �verf�ra inst�llningar fr�n MTCP.CFG till WATTCP.CFG.
Keywords:    mTCP, WATTCP, DHCP
End
