Begin3
Language:    SV, 850, Swedish
Title:       CTMouse
Description: FreeDOS musdrivrutin
Keywords:    Mus, hjul
End
