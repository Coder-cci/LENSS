Begin3
Language:    SV, 850, Swedish
Title:       fc
Description: Filj�mf�relseverktyg
Keywords:    freedos, fil, j�mf�relse, fc
End
