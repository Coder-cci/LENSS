Begin3
Language:    SV, 850, Swedish
Title:       sleep
Description: sleep liknar UNIX-verktyget med samma namn. sleep kan anv�ndas f�r att pausa k�rningen av kommandofiler en studn. sleep ger tillbaka tid till operativsystem som har st�d f�r det. sleep k�nner igen och respekterar DOS switchar.
Keywords:    ut�kning, verktyg, f�rdr�jning
End
