Begin3
Language:    SV, 850, Swedish
Title:       cURL
Description: Curl �r ett kommandoradsverktyg f�r att �verf�ra data angiven med URL-syntax.
Keywords:    freedos, curl
End
