Begin3
Language:    SV, 850, Swedish
Title:       FreeCom
Description: FreeDOS kommandoskal
Keywords:    freecom freedos kommandoskal
End
