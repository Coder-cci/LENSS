Begin3
Language:    SV, 850, Swedish
Title:       Mirror Magic
Description: Ett spel i arkadstil likt Deflektor (C 64) eller Mindbender (Amiga)
End
