Begin3
Language:    SV, 850, Swedish
Title:       sort
Description: Sortera inneh�llet i en textfil, sortera valfritt enligt NLS-tabell 
Keywords:    sorter, text, fil
End
