vchkbox [flaggor]

   tba         (Fortfarande under utveckling, mer kommer att annonseras)
