Begin3
Language:    SV, 850, Swedish
Title:       KEYB layouter
Description: Tangentbordslayouter f�r KEYB
Keywords:    keyb,layouter
End
