Begin3
Language:    SV, 850, Swedish
Title:       attrib
Description: Visa och s�tt filattribut
Keywords:    freedos, attrib
End
