FDSHELL

FDSHELL �r en �ppenk�llkodsversion av Microsofts grafiska anv�ndargr�nssnitt DOSSHELL
Modifiera DOSSHELL.INI om det beh�vs

