Begin3
Language:    SV, 850, Swedish
Title:       HIMEMSX
Description: HimemSX �r en gren av HimemX. Dess huvudfunktion �r att den kan hantera mer �n 4 Gbyte minne.
Keywords:    ut�kat minne, himem, himemsx, minneshanterarer, superut�kat, XMS
End
