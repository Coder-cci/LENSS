Begin3
Language:    SV, 850, Swedish
Title:       RDISK
Description: RDISK �r en drivrutin som skapar en RAM-disk av upp till 2GB XMS-minne.
Keywords:    disk, drivrutin, minne, ramdisk, rdisk, xms
End
