Begin3
Language:    SV, 850, Swedish
Title:       SSH2DOS
Description: SSH-klient f�r SSH-protokoll version 2.0. Inneh�ller ocks� SCP, SFTP och telnet i b�de 8086- och 386-versioner.
Keywords:    ssh protokoll n�tverk kommunikation fj�rr�tkomst
End
