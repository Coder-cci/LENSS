Begin3
Language:    SV, 850, Swedish
Title:       LAME
Description: Verktyg f�r att manipulera MP3-musikfiler, inklusive konvertering till andra format och dekomprimering till .WAV.
Keywords:    mp3, lame, konvertera, ljud, wav
End
