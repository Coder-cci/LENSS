Begin3
Language:    SV, 850, Swedish
Title:       Links
Description: Links �r en Lynx-liknande text och grafisk WWW-l�sare.
Keywords:    www, l�sare, internet
End
