Begin3
Language:    SV, 850, Swedish
Title:       ping
Description: Verktyget ping f�r internetdiagnostik. Denna version extraherades fr�n Watt-32 v2.2-sviten.
Keywords:    ping
End
