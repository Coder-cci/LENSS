Begin3
Language:    SV, 850, Swedish
Title:       FreeDOS-hj�lp (AMB)
Description: FreeDOS-hj�lpfiler i AMB -ormat
Keywords:    freedos, hj�lp, dokument, text, amb
End
