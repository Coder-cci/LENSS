Begin3
Language:    SV, 850, Swedish
Title:       Uptime (Chamorro)
Description: Rapporterar k�rtid, �ven inuti DOSEmu. Liknar uptime i UNIX.
Summary:     UPTIME �r ett 16-bitars DOS-verktyg som visar systems k�rtid genom att automatiskt detektera n�r det f�rst startades. Det duplicerar *NIX uptime, en av de mest grundl�ggande UNIX-kommandona vilket l�ter dig snabbt bekr�fta hur l�nge ditt system har varit upp och k�rt sedan det senast startade eller startades om.
Keywords:    k�rtid
End
