Begin3
Language:    SV, 850, Swedish
Title:       Lzip
Description: En datakomprimerare baserad p� LZMS-algoritmen.
Keywords:    kommando.com, skal, interaktivt
End
