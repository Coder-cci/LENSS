Begin3
Language:    SV, 850, Swedish
Title:       BZIP2
Description: BZIP2-kompressionprogram
Keywords:    bzip, bunzip, zip, unzip, komprimerare
End
