vinsert [flaggor]

Infoga en tomrad p� aktuell position.

    [inga]      Infoga en tom rad.
    n           Infoga n tomma rader.
    /A n        S�tt textattribut till n.
    /B f�rg     S�tt textattribut f�r bakgrunden till f�rg (eller v�rde).
    /F f�rg     S�tt textattribut f�r f�rgrunden till f�rg (eller v�rde).
    /G          Global infogning.
    /L          Lokal infogning. (Standard)
    /K n        Anv�nd n ist�llet f�r ramtecken f�r att identifiera ramar.

