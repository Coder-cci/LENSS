Begin3
Language:    SV, 850, Swedish
Title:       JEMM386
Description: Jemm386 �r en expanderad minneshanterare f�r DOS
Summary:     Jemm386 �r en expanderad minneshanterare f�r DOS, baserad p� k�llkoden f�r FreeDOS EMM386. Den har flera f�rdelar j�mf�r med EMM386 fr�n FreeDOS och/eller MS-DOS. Den beh�ver endast 192 byte DOS-minne, den beh�ver v�ldig lite ut�kat minne, den �r snabbare, den fugnerar med MS-DOS, FreeDOS och EDR-DOS, den anv�nder funktioner implementerade i senare CPU:er f�r att f�rb�ttr prestanda, till skillnad fr�n FreeDOS Emm386 har Jemm386 fullst�ndigt VDS-st�d, den kan l�sas in fr�n kommandoraden.
Keywords:    HIMEM + EMM386, STABIL, KOMPATIBILITET, minneshanterare, jemmex, himemx
End
