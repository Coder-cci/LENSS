Begin3
Language:    SV, 850, Swedish
Title:       7-ZIP
Description: p7zip �r en snabb portering av 7za.exe (kommandoradsversionen av 7zip). 7-Zip �r ett filarkveringsprogram med den h�gsta kompressiongraden.
Keywords:    7zip, p7zip, komprimering, zip, unzip, arj
End
