Begin3
Language:    SV, 850, Swedish
Title:       Senet
Description: Ett mycket gamalt spel som daterar tillbaka till forntida Egypten
Summary:     Senet �r ett mycket gamlat spel, som g�r tillbaka till det gamla Egypten. Eftersom det �r s� gamalt och ingen i forntida Egypten bevarade reglerna �t senare generationer �r de exakta reglerna n�got av ett mysterium. Historiker har f�rs�kt lista ut reglerna i Senet, men de �r oense om detaljerna.
Keywords:    Spel
End
