Begin3
Language:    SV, 850, Swedish
Title:       LABEL
Description: S�tter eller �ndrar diskens volymetikett
Keywords:    etikett, diskvolym
End
