Begin3
Language:    SV, 850, Swedish
Title:       zoo
Description: Manipulera zoo-arkiv.
Keywords:    zoo
End
