Begin3
Language:    SV, 850, Swedish
Title:       USBDOS
Description: Samling DOS-drivrutiner f�r UHCI (USB 1.1 12Mbit/1.5Mbit)
Keywords:    DOS USB drivrutin tangentbord musport uhci ohci ehci xhci
End
