Begin3
Language:    SV, 850, Swedish
Description: S�tter DOS-versionen under ett programs k�rning.
End
