Begin3
Language:    SV, 850, Swedish
Title:       WATTCP
Description: WATTCP
Keywords:    freedos, curl
End
