Begin3
Language:    SV, 850, Swedish
Title:       Liquid War
Description: Ett unikt krigsspel f�r flera spelare.
End
