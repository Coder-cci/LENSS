Begin3
Language:    SV, 850, Swedish
Title:       Defrag
Description: Defragmenteringsverktyg.
Keywords:    defragmenterare
End
