Begin3
Language:    SV, 850, Swedish
Title:       Iter Vehems ad Necem
Description: Ett grafiskt rogue-liknande spel.
End
