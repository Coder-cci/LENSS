Begin3
Language:    SV, 850, Swedish
Title:       DOSMid
Description: MIDI-spelare f�r m�nga synthesizrar (AWE, MPU-401, OPL...)
Summary:     DOSMid �r en MIDI- och MUS-spelare f�r DOS. Det �r en real mode-applikation designad f�r att k�ra p� mycket sm� h�rdvarukonfigurationer. Den spelar standard MIDI-filer s� v�l som MIDI i RIFF (d.v.s RMID) och MUS-l�tar (anv�nda av Id Software i flertalet spel, t.ex. Doom, Heretic, Hexen o.s.v.).
Keywords:    midi,mus,rmid,spelare
End
