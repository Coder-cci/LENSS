Begin3
Language:    SV, 850, Swedish
Title:       FreeDOS hj�lpprogram
Description: Kommandofiler f�r att utf�ra diverse uppgifter i FreeDOS
Summary:     Kommandofiler som utf�r uppgifter. I stil med meddelandet 'V�lkommen till FreeDOS', CD/DVD-ROM-initiering med mera
Keywords:    uppstart cd dvd spr�k meddelanden autoexec config system drivrutin ut�kning
End
