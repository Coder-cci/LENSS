Begin3
Language:    SV, 850, Swedish
Title:       Bolitaire
Description: En DOS-klon av Freecel 
End
