# edlin.sv - Swedish-language messages file
#
# Author: Gregory Pietsch
#
# DESCRIPTION:
#
# This file contains #defines for all the message strings in edlin.
# For internationalization fun, just translate the messages in this
# file.
# Swedish translation Oct 2006 /A.J
# Updated translation Dec 2021 /Sebastian Rasmussen

1.0:Jj
1.1::\040:\040
1.2:OK?\040
1.3:Inmatningsfil
1.4:%s: %lu rad inl�st\n
1.5:%s: %lu rader inl�sta\n
1.6:%s: %lu rad skriven\n
1.7:%s: %lu rader skrivna\n
1.8:%lu:%c%s\n
1.9:Tryck <retur> 
1.10:%lu:\040
1.11:Hittades ej
1.12:%lu: %s\n
1.13:\nedlin har f�ljande kommandon:\n
1.14:#                 redigera en rad       [#],[#],#m        flytta
1.15:a                 l�gg till p� slutet   [#][,#]p          sida
1.16:[#],[#],#,[#]c    kopiera               q                 avsluta
1.17:[#][,#]d          ta bort               [#][,#][?]r$,$    ers�tt
1.18:e<>               avsluta (spara)       [#][,#][?]s$      s�k
1.19:[#]i              infoga                [#]t<>            �verf�r
1.20:[#][,#]l          lista                 [#]w<>            spara\n
1.21:d�r $ �r en str�ng, <> �r ett filnamn,
1.22:# �r ett radnummer (.=aktuell rad, $=sista raden,
1.23: uttryck med +/- kan anv�ndas)\n
1.24:, copyright (c) 2003 Gregory Pietsch
1.25:Detta program kommer utan N�GON SOM HELST GARANTI.
1.26:Det h�r �r fri programvara, och du f�r g�rna distribuera
1.27:det vidare under villkoren f�r GNU General Public License
1.28:antingen version 2 av licensen, eller om du vill n�gon senare
1.29:version.\n
1.30:Slut p� minne
1.31:Felaktig str�ngl�ngd
1.32:Felaktig str�ngposition
1.33:F�rst�r ej, skriv ? f�r hj�lp.
1.34:Filnamn saknas
1.35:F�r stor buffert
1.36:Ogiltig buffertposition
1.37:FEL: %s\n

# END OF FILE
