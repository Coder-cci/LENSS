Begin3
Language:    SV, 850, Swedish
Title:       DOS Defender
Description: DOS Defender �r ett x86 Real Mode-spel f�r DOS f�r Ludum Dare #31 (December, 2014). Eftersom endas ett f�tal DOS-maskiner fortfarande existerar �r m�lplattformen egentligen DOSBox, men det b�r fungera i viss utstr�ckning p� vilket DOS-system som helst. Spelet kan spelas med musen men �r avsett att spelas med en joystick/spelkontroll.
Keywords:    spel
End
