Begin3
Language:    SV, 850, Swedish
Title:       LZMA-verktyg
Description: Arbetar med .lzma-komprimerade filer (skiljer sig fr�n 7-zip)
Keywords:    lzma
End
