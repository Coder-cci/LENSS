Begin3
Language:    SV, 850, Swedish
Title:       Tree
Description: Visar katalogstrukturen grafiskt f�r en enhet eller s�kv�g.
Summary:     Visar grafiskt mappstrukturen f�r en enhet eller s�kv�g. St�d f�r meddelandekataloger (olika spr�k) via cats och kan kompileras f�r b�de Windows NT/9x och DOS.
Keywords:    tr�d, FreeDOS, DOS, Win32
End
