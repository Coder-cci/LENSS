vmath [flaggor]

Super enkelt matteverktyg. Det �r INTE en kalkylator och �r begr�nsat till att
arbeta p� tal mellan 0-32767. Bra f�r loopar, best�mma sk�rmpositioner etc.

    +, ADD      L�gg till n�sta nummer till summan.
    -, SUB      Subtrahera n�sta nummer fr�n summan.
    *, MUL      Multiplicera summa med n�sta nummer.
    /, DIV      Dividera summa med n�sta nummer.
    \, MOD      Dividera summa med n�sta nummer och s�tt summan till resten.
    AND         Logiskt OCH.
    OR          Logiskt ELLER.
    XOR         Logiskt exklusivt ELLER.
    SHR         Bitskiftning �t h�ger
    SHL         Bitskiftning �t v�nster.

    /H          S�tt utmatning till hexadecimalt.
    /D          S�tt utmatning till decimalt.
