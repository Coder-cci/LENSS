Begin3
Language:    SV, 850, Swedish
Description: En fullt konfigurerbar programstartare med flera menyer f�r DOS. Det inkluderar ocks� Font Designer och flera andra verktyg. (Kr�ver mus)
Keywords:    dos starta program efntdsgn meny kiosk 16-bit
End
