Begin3
Language:    SV, 850, Swedish
Title:       FDAPM
Description: APM/ACPI styrning/info, str�mspar TSR/styrning, cachet�mning, omstart... {en ers�ttare f�r MS-DOS POWER}
Keywords:    APM, ACPI, str�m, batteri, str�mspar, spinna ner, dpms-sk�rm, begr�nsa hastighet, starta om, st�ng ner
End
