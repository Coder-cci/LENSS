Begin3
Language:    SV, 850, Swedish
Title:       DISPLAY
Description: FreeDOS drivrutin f�r kodsideshantering (sk�rm eller skrivare)
Keywords:    visa, ega, vga, nls, cpi, cpx
End
