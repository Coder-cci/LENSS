Begin3
Language:    SV, 850, Swedish
Title:       cal
Description: Kalenderprogram, i stil med UNIX cal
Keywords:    freedos
End
