Begin3
Language:    SV, 850, Swedish
Title:       Vertigo
Description: Flygsimulator som fokuserar p� realism i flygmodellen.
End
