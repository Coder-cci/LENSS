Begin3
Language:    SV, 850, Swedish
Title:       DEBUG
Description: Ett verktyg f�r programtestning och redigering
Keywords:    32-bitars avlusare, fels�kning, avlusare, DPMI-avlusare, k�rnavlusare
End
