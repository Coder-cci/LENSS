Begin3
Language:    SV, 850, Swedish
Title:       mode
Description: S�tt l�get f�r dina enheter:
Summary:     S�tt l�get f�r dina enheter:|- skicka ESC/P kontrollkoder f�r 80/132-kolumner och 6/8-rader per tum till skrivare|- omdirigera skrivare till NUL eller serieport|- s�tt serieportsparametrar|- g�r kodsides�tg�rder och visa DISPLAY-status|- v�lj 40/80/132x25/28/43/50/60-sk�rml�ge eller v�lj x8/14/16-typsnitt, tillg�nglighet beroende p� din|h�rdvara. Skifta CGA-sk�rmen sidledes.|- styr och kontrollera switchar och l�sstatus p� tangentbordet (num/...)|- styr tangentbordets repetitionshastighet och f�rdr�jning
Keywords:    freedos, mode, l�ge, visa
End
