Begin3
Language:    SV, 850, Swedish
Title:       SAMCFG
Description: En upps�ttning av exempelfiler f�r att skapa C:CONFIG.SYS och C:AUTOEXEC.BAT
Keywords:    freedos, exempel, konfiguration, config.sys, autoexec.bat, kommandofil, skript
End
