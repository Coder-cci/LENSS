Begin3
Language:    SV, 850, Swedish
Title:       Arachne
Description: en webbl�sare f�r DOS (8086- & i386-versioner)
Keywords:    n�tverk, www, webbl�sare
End
