Begin3
Language:    SV, 850, Swedish
Title:       GNU grep
Description: grep genoms�ker filer (eller standard in) efter rader som matcar ett givet m�nster. M�nstret kan vara ett regulj�rt uttryck eller en bokstavlig str�ng.
Keywords:    grep,m�nster
End
