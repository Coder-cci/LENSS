Begin3
Language:    SV, 850, Swedish
Title:       FreeDOS hj�lp (HTML)
Description: HTML-visare och inneh�ll f�r FreeDOS-hj�lp
Keywords:    hj�lp, html
End
