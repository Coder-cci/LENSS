Begin3
Language:    SV, 850, Swedish
Title:       DU
Description: Visa diskanv�ndning, i stil med du under UNIX
Keywords:    du, visa diskanv�ndning
End
