Begin3
Language:    SV, 850, Swedish
Title:       E100PKT
Description: Paketdrivrutin f�r DOS
Keywords:    n�tverk, ethernet, paket, drivrutin, e100, intel
End
