Begin3
Language:    SV, 850, Swedish
Title:       swsubst
Description: SUBST och JOIN
Keywords:    freedos, subst, join
End
