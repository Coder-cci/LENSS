Begin3
Language:    SV, 850, Swedish
Title:       TEE
Description: Sparar en kopia av dess indata till en fil, medan en kopia skrivs ut p� stdout
Keywords:    tee, unix
End
