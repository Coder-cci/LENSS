Begin3
Language:    SV, 850, Swedish
Description: DOS Navigator 2 �ppen k�llkod�r en filhanterare baserad p� DOS Navigator (c) 1991-99 av RIT Research Labs.
End
