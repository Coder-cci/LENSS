Begin3
Language:    SV, 850, Swedish
Title:       mTCP (upx)
Description: En UPX:ad samling TCP/IP-verktyg f�r 16-bitars DOS: DHCP, IRC, FTP, Telnet, Netcat, HTGet, Ping, SNTP
Keywords:    dos tcp/ip realmode dhcp ftp telnet htget irc ircjr netcat sntp ping �ppen k�llkod 16-bitars
End
