Begin3
Language:    SV, 850, Swedish
Title:       Lynx
Description: Lynx text och grafik WWW-l�sare (DJGPP-portering)
Summary:     Lynx WWW-l�sare f�r text- och grafikl�ge (DJGPP-portering, inkluderar noise v0.6.3-beta)
Keywords:    www, l�sare, internet
End
