Begin3
Language:    SV, 850, Swedish
Title:       HTGET
Description: HTGET �r en filh�mtare som h�mtar filer fr�n HTTP-servrar.
Keywords:    freedos, htget
End
