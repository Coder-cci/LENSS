Begin3
Language:    SV, 850, Swedish
Title:       E1000PKT
Description: Paketdrivrutin f�r Intel(R) PRO/1000-kort, t.ex. 82544-, 82540-, 82545-, 82541- och 82547-baserade Ethernet kontrollerkort.
Keywords:    82544, 82540, 82545, 82541, 82547, GIGPKTDRVR, Gigabit paketdrivrutin
End
