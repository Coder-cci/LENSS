Begin3
Language:    SV, 850, Swedish
Title:       Format
Description: Diskformateringsprogram -- skapar FAT-filsystem och l�gniv�formaterar disketter
Keywords:    freedos, format, fat12, fat16, fat32, diskett, h�rddisk, spegling, oformatera
End
