# Hj�lpmeddelanden

0.0:Move
0.1:Flytter en fil/katalog till en annan plats.
0.2:(C) 1997-2002 by Joe Cosentino
0.3:(C) 2003-2004 by Imre Leber
0.4:Syntax: MOVE
0.5:k�lla1[, k�lla2[,...]] destination
0.6: k�lla       Namnet p� filen eller katalogen du vill flytta (byta namn p�)
0.7: destination Vart du vill flytta filen/filerna
0.8:          Undertrycker f�rfr�gan om du vill skriva �ver
0.9:             en existerande destinations fil.
0.10:         Ser till att f�rfr�gan sker om �verskrivning av
0.11:             existerande destinationsfil.
0.12:          Verifierar varje file d� den skrivs till destinationsfilen
0.13:             f�r att s�kerst�lla att destinations filerna �r identiska med
0.14:             k�llfilerna
0.15:Not:
0.16:Du kan flytta kataloger med detta verktyg

# Diverse meddelanden

1.0:finns ej!
1.1:finns redan!
1.2:Skriv �ver fil
1.3:Problem vid f�rflyttning av katalog
1.4:Problem vid f�rflyttning av fil
1.5:Ogiltig parameter
1.6:Ogiltig enhetsspecifikation f�r k�lla
1.7:Ogiltig destinationsfil
1.8: finns inte som en katalog. Skapa den?
1.9:Ogiltig k�llfil
1.10:Kan inte skapa katalog
1.11:Fil kan inte kopieras ovanp� sig sj�lv
1.12:Kan inte flytta en fil till en katalog
1.13:Fil finns redan
1.14:Fil kan inte kopieras ovanp� sig sj�lv
1.15:�tkomst nekad
1.16:Otillr�ckligt diskutrymme i destinationss�kv�g
1.17:Otillr�ckligt diskutrymme
1.18:N�dv�ndig parameter saknas
1.19:Ogiltig k�llspecifikation
1.20:K�lls�kv�g finns inte
1.21:K�lls�kv�g f�r l�ng\n
1.22:Destinationss�kv�g f�r l�ng\n
1.23:Ogiltig enhetsspecifikation f�r destination\n
1.24:Destinationss�kv�g f�r l�ng\n
1.25:Kan inte �ppna k�llfil
1.26:Kan inte skapa destinationsfil
1.27:Skrivfel vid destinationsfil
1.28:Kan inte skapa katalog
1.29:Otillr�ckligt diskutrymme i destinationss�kv�g

# J/N/Alla/Inga; Enkla meddelanden

2.0:J
2.1:N
2.2:Alla
2.3:Inga
2.4:ok
