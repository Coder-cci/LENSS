Begin3
Language:    SV, 850, Swedish
Title:       UNFORMAT
Description: Unformat kan �terst�lla en disk som du formaterat av misstag.
Keywords:    format, unformat, h�rddisk,
End
