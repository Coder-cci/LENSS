vver [flaggor]

V8Power informationsprogram.

    [inga]      Skriver ut all information till STDOUT.
    all         Skriver ut all information till STDOUT.
    title       Skriver ut fullst�ndig titel till STDOUT.
    copyright   Skriver ut upphovsr�ttsmeddelande till STDOUT.
    version     Skriver ut versionsinformation till STDOUT.
    license     Skriver ut licensinformation till STDOUT.
    url         Skriver ut url till webbplats till STDOUT.
    email       Skriver ut e-postadress till STDOUT.
