Begin3
Language:    SV, 850, Swedish
Title:       Smiley
Description: Ett enkelt spel i pong-stil (VGA, 386+)
Summary:     Ett enkelt spel i pong-stil mestadels f�r att testa olika aspected av Danger Engine. Kr�ver VGA och 386+. En mus rekommenderas starkt.
Keywords:    dos spel
End
