Begin3
Language:    SV, 850, Swedish
Title:       ElTorito
Description: Enkelt paket f�r SysLinux ElToritor CD-drivrutin.
End
