Begin3
Language:    SV, 850, Swedish
Title:       RECOVER
Description: �terst�ller diskar eller f�rlorad filer.
Keywords:    �terst�ll, diskar, filer
End
