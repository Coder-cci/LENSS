Begin3
Language:    SV, 850, Swedish
Title:       terminal
Description: En liten vt100/ansi-terminale f�r varje pc
Keywords:    terminal, rs-232, vt100
End
